

module ADC(input RES_HARD, input CLK, input CS, input LOCK, input CONVECT, input BYTESWAP
			  output BYSY, output [7 : 0]DATA );
			  
			  
			  
endmodule			  